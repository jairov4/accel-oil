library verilog;
use verilog.vl_types.all;
entity nfa_accept_samples_generic_hw_top is
    generic(
        C_nfa_initials_buckets_REMOTE_DESTINATION_ADDRESS: integer := 0;
        C_nfa_initials_buckets_AWIDTH: integer := 32;
        C_nfa_initials_buckets_DWIDTH: integer := 64;
        C_nfa_initials_buckets_NATIVE_DWIDTH: integer := 64;
        C_nfa_finals_buckets_REMOTE_DESTINATION_ADDRESS: integer := 0;
        C_nfa_finals_buckets_AWIDTH: integer := 32;
        C_nfa_finals_buckets_DWIDTH: integer := 64;
        C_nfa_finals_buckets_NATIVE_DWIDTH: integer := 64;
        C_nfa_forward_buckets_REMOTE_DESTINATION_ADDRESS: integer := 0;
        C_nfa_forward_buckets_AWIDTH: integer := 32;
        C_nfa_forward_buckets_DWIDTH: integer := 64;
        C_nfa_forward_buckets_NATIVE_DWIDTH: integer := 64;
        C_sample_buffer_REMOTE_DESTINATION_ADDRESS: integer := 0;
        C_sample_buffer_AWIDTH: integer := 32;
        C_sample_buffer_DWIDTH: integer := 64;
        C_sample_buffer_NATIVE_DWIDTH: integer := 64;
        C_indices_REMOTE_DESTINATION_ADDRESS: integer := 0;
        C_indices_AWIDTH: integer := 32;
        C_indices_DWIDTH: integer := 64;
        C_indices_NATIVE_DWIDTH: integer := 64;
        C_SPLB_SLV0_BASEADDR: integer := 0;
        C_SPLB_SLV0_HIGHADDR: integer := 15;
        C_SPLB_SLV0_AWIDTH: integer := 32;
        C_SPLB_SLV0_DWIDTH: integer := 32;
        C_SPLB_SLV0_NUM_MASTERS: integer := 8;
        C_SPLB_SLV0_MID_WIDTH: integer := 3;
        C_SPLB_SLV0_NATIVE_DWIDTH: integer := 32;
        C_SPLB_SLV0_P2P : integer := 0;
        C_SPLB_SLV0_SUPPORT_BURSTS: integer := 0;
        C_SPLB_SLV0_SMALLEST_MASTER: integer := 32;
        C_SPLB_SLV0_INCLUDE_DPHASE_TIMER: integer := 0;
        RESET_ACTIVE_LOW: integer := 1
    );
    port(
        nfa_initials_buckets_MPLB_Clk: in     vl_logic;
        nfa_initials_buckets_MPLB_Rst: in     vl_logic;
        nfa_initials_buckets_M_request: out    vl_logic;
        nfa_initials_buckets_M_priority: out    vl_logic_vector(1 downto 0);
        nfa_initials_buckets_M_busLock: out    vl_logic;
        nfa_initials_buckets_M_RNW: out    vl_logic;
        nfa_initials_buckets_M_BE: out    vl_logic_vector;
        nfa_initials_buckets_M_MSize: out    vl_logic_vector(1 downto 0);
        nfa_initials_buckets_M_size: out    vl_logic_vector(3 downto 0);
        nfa_initials_buckets_M_type: out    vl_logic_vector(2 downto 0);
        nfa_initials_buckets_M_TAttribute: out    vl_logic_vector(15 downto 0);
        nfa_initials_buckets_M_lockErr: out    vl_logic;
        nfa_initials_buckets_M_abort: out    vl_logic;
        nfa_initials_buckets_M_UABus: out    vl_logic_vector(31 downto 0);
        nfa_initials_buckets_M_ABus: out    vl_logic_vector(31 downto 0);
        nfa_initials_buckets_M_wrDBus: out    vl_logic_vector;
        nfa_initials_buckets_M_wrBurst: out    vl_logic;
        nfa_initials_buckets_M_rdBurst: out    vl_logic;
        nfa_initials_buckets_PLB_MAddrAck: in     vl_logic;
        nfa_initials_buckets_PLB_MSSize: in     vl_logic_vector(1 downto 0);
        nfa_initials_buckets_PLB_MRearbitrate: in     vl_logic;
        nfa_initials_buckets_PLB_MTimeout: in     vl_logic;
        nfa_initials_buckets_PLB_MBusy: in     vl_logic;
        nfa_initials_buckets_PLB_MRdErr: in     vl_logic;
        nfa_initials_buckets_PLB_MWrErr: in     vl_logic;
        nfa_initials_buckets_PLB_MIRQ: in     vl_logic;
        nfa_initials_buckets_PLB_MRdDBus: in     vl_logic_vector;
        nfa_initials_buckets_PLB_MRdWdAddr: in     vl_logic_vector(3 downto 0);
        nfa_initials_buckets_PLB_MRdDAck: in     vl_logic;
        nfa_initials_buckets_PLB_MRdBTerm: in     vl_logic;
        nfa_initials_buckets_PLB_MWrDAck: in     vl_logic;
        nfa_initials_buckets_PLB_MWrBTerm: in     vl_logic;
        nfa_finals_buckets_MPLB_Clk: in     vl_logic;
        nfa_finals_buckets_MPLB_Rst: in     vl_logic;
        nfa_finals_buckets_M_request: out    vl_logic;
        nfa_finals_buckets_M_priority: out    vl_logic_vector(1 downto 0);
        nfa_finals_buckets_M_busLock: out    vl_logic;
        nfa_finals_buckets_M_RNW: out    vl_logic;
        nfa_finals_buckets_M_BE: out    vl_logic_vector;
        nfa_finals_buckets_M_MSize: out    vl_logic_vector(1 downto 0);
        nfa_finals_buckets_M_size: out    vl_logic_vector(3 downto 0);
        nfa_finals_buckets_M_type: out    vl_logic_vector(2 downto 0);
        nfa_finals_buckets_M_TAttribute: out    vl_logic_vector(15 downto 0);
        nfa_finals_buckets_M_lockErr: out    vl_logic;
        nfa_finals_buckets_M_abort: out    vl_logic;
        nfa_finals_buckets_M_UABus: out    vl_logic_vector(31 downto 0);
        nfa_finals_buckets_M_ABus: out    vl_logic_vector(31 downto 0);
        nfa_finals_buckets_M_wrDBus: out    vl_logic_vector;
        nfa_finals_buckets_M_wrBurst: out    vl_logic;
        nfa_finals_buckets_M_rdBurst: out    vl_logic;
        nfa_finals_buckets_PLB_MAddrAck: in     vl_logic;
        nfa_finals_buckets_PLB_MSSize: in     vl_logic_vector(1 downto 0);
        nfa_finals_buckets_PLB_MRearbitrate: in     vl_logic;
        nfa_finals_buckets_PLB_MTimeout: in     vl_logic;
        nfa_finals_buckets_PLB_MBusy: in     vl_logic;
        nfa_finals_buckets_PLB_MRdErr: in     vl_logic;
        nfa_finals_buckets_PLB_MWrErr: in     vl_logic;
        nfa_finals_buckets_PLB_MIRQ: in     vl_logic;
        nfa_finals_buckets_PLB_MRdDBus: in     vl_logic_vector;
        nfa_finals_buckets_PLB_MRdWdAddr: in     vl_logic_vector(3 downto 0);
        nfa_finals_buckets_PLB_MRdDAck: in     vl_logic;
        nfa_finals_buckets_PLB_MRdBTerm: in     vl_logic;
        nfa_finals_buckets_PLB_MWrDAck: in     vl_logic;
        nfa_finals_buckets_PLB_MWrBTerm: in     vl_logic;
        nfa_forward_buckets_MPLB_Clk: in     vl_logic;
        nfa_forward_buckets_MPLB_Rst: in     vl_logic;
        nfa_forward_buckets_M_request: out    vl_logic;
        nfa_forward_buckets_M_priority: out    vl_logic_vector(1 downto 0);
        nfa_forward_buckets_M_busLock: out    vl_logic;
        nfa_forward_buckets_M_RNW: out    vl_logic;
        nfa_forward_buckets_M_BE: out    vl_logic_vector;
        nfa_forward_buckets_M_MSize: out    vl_logic_vector(1 downto 0);
        nfa_forward_buckets_M_size: out    vl_logic_vector(3 downto 0);
        nfa_forward_buckets_M_type: out    vl_logic_vector(2 downto 0);
        nfa_forward_buckets_M_TAttribute: out    vl_logic_vector(15 downto 0);
        nfa_forward_buckets_M_lockErr: out    vl_logic;
        nfa_forward_buckets_M_abort: out    vl_logic;
        nfa_forward_buckets_M_UABus: out    vl_logic_vector(31 downto 0);
        nfa_forward_buckets_M_ABus: out    vl_logic_vector(31 downto 0);
        nfa_forward_buckets_M_wrDBus: out    vl_logic_vector;
        nfa_forward_buckets_M_wrBurst: out    vl_logic;
        nfa_forward_buckets_M_rdBurst: out    vl_logic;
        nfa_forward_buckets_PLB_MAddrAck: in     vl_logic;
        nfa_forward_buckets_PLB_MSSize: in     vl_logic_vector(1 downto 0);
        nfa_forward_buckets_PLB_MRearbitrate: in     vl_logic;
        nfa_forward_buckets_PLB_MTimeout: in     vl_logic;
        nfa_forward_buckets_PLB_MBusy: in     vl_logic;
        nfa_forward_buckets_PLB_MRdErr: in     vl_logic;
        nfa_forward_buckets_PLB_MWrErr: in     vl_logic;
        nfa_forward_buckets_PLB_MIRQ: in     vl_logic;
        nfa_forward_buckets_PLB_MRdDBus: in     vl_logic_vector;
        nfa_forward_buckets_PLB_MRdWdAddr: in     vl_logic_vector(3 downto 0);
        nfa_forward_buckets_PLB_MRdDAck: in     vl_logic;
        nfa_forward_buckets_PLB_MRdBTerm: in     vl_logic;
        nfa_forward_buckets_PLB_MWrDAck: in     vl_logic;
        nfa_forward_buckets_PLB_MWrBTerm: in     vl_logic;
        sample_buffer_MPLB_Clk: in     vl_logic;
        sample_buffer_MPLB_Rst: in     vl_logic;
        sample_buffer_M_request: out    vl_logic;
        sample_buffer_M_priority: out    vl_logic_vector(1 downto 0);
        sample_buffer_M_busLock: out    vl_logic;
        sample_buffer_M_RNW: out    vl_logic;
        sample_buffer_M_BE: out    vl_logic_vector;
        sample_buffer_M_MSize: out    vl_logic_vector(1 downto 0);
        sample_buffer_M_size: out    vl_logic_vector(3 downto 0);
        sample_buffer_M_type: out    vl_logic_vector(2 downto 0);
        sample_buffer_M_TAttribute: out    vl_logic_vector(15 downto 0);
        sample_buffer_M_lockErr: out    vl_logic;
        sample_buffer_M_abort: out    vl_logic;
        sample_buffer_M_UABus: out    vl_logic_vector(31 downto 0);
        sample_buffer_M_ABus: out    vl_logic_vector(31 downto 0);
        sample_buffer_M_wrDBus: out    vl_logic_vector;
        sample_buffer_M_wrBurst: out    vl_logic;
        sample_buffer_M_rdBurst: out    vl_logic;
        sample_buffer_PLB_MAddrAck: in     vl_logic;
        sample_buffer_PLB_MSSize: in     vl_logic_vector(1 downto 0);
        sample_buffer_PLB_MRearbitrate: in     vl_logic;
        sample_buffer_PLB_MTimeout: in     vl_logic;
        sample_buffer_PLB_MBusy: in     vl_logic;
        sample_buffer_PLB_MRdErr: in     vl_logic;
        sample_buffer_PLB_MWrErr: in     vl_logic;
        sample_buffer_PLB_MIRQ: in     vl_logic;
        sample_buffer_PLB_MRdDBus: in     vl_logic_vector;
        sample_buffer_PLB_MRdWdAddr: in     vl_logic_vector(3 downto 0);
        sample_buffer_PLB_MRdDAck: in     vl_logic;
        sample_buffer_PLB_MRdBTerm: in     vl_logic;
        sample_buffer_PLB_MWrDAck: in     vl_logic;
        sample_buffer_PLB_MWrBTerm: in     vl_logic;
        indices_MPLB_Clk: in     vl_logic;
        indices_MPLB_Rst: in     vl_logic;
        indices_M_request: out    vl_logic;
        indices_M_priority: out    vl_logic_vector(1 downto 0);
        indices_M_busLock: out    vl_logic;
        indices_M_RNW   : out    vl_logic;
        indices_M_BE    : out    vl_logic_vector;
        indices_M_MSize : out    vl_logic_vector(1 downto 0);
        indices_M_size  : out    vl_logic_vector(3 downto 0);
        indices_M_type  : out    vl_logic_vector(2 downto 0);
        indices_M_TAttribute: out    vl_logic_vector(15 downto 0);
        indices_M_lockErr: out    vl_logic;
        indices_M_abort : out    vl_logic;
        indices_M_UABus : out    vl_logic_vector(31 downto 0);
        indices_M_ABus  : out    vl_logic_vector(31 downto 0);
        indices_M_wrDBus: out    vl_logic_vector;
        indices_M_wrBurst: out    vl_logic;
        indices_M_rdBurst: out    vl_logic;
        indices_PLB_MAddrAck: in     vl_logic;
        indices_PLB_MSSize: in     vl_logic_vector(1 downto 0);
        indices_PLB_MRearbitrate: in     vl_logic;
        indices_PLB_MTimeout: in     vl_logic;
        indices_PLB_MBusy: in     vl_logic;
        indices_PLB_MRdErr: in     vl_logic;
        indices_PLB_MWrErr: in     vl_logic;
        indices_PLB_MIRQ: in     vl_logic;
        indices_PLB_MRdDBus: in     vl_logic_vector;
        indices_PLB_MRdWdAddr: in     vl_logic_vector(3 downto 0);
        indices_PLB_MRdDAck: in     vl_logic;
        indices_PLB_MRdBTerm: in     vl_logic;
        indices_PLB_MWrDAck: in     vl_logic;
        indices_PLB_MWrBTerm: in     vl_logic;
        splb_slv0_SPLB_Clk: in     vl_logic;
        splb_slv0_SPLB_Rst: in     vl_logic;
        splb_slv0_PLB_ABus: in     vl_logic_vector(31 downto 0);
        splb_slv0_PLB_UABus: in     vl_logic_vector(31 downto 0);
        splb_slv0_PLB_PAValid: in     vl_logic;
        splb_slv0_PLB_SAValid: in     vl_logic;
        splb_slv0_PLB_rdPrim: in     vl_logic;
        splb_slv0_PLB_wrPrim: in     vl_logic;
        splb_slv0_PLB_masterID: in     vl_logic_vector;
        splb_slv0_PLB_abort: in     vl_logic;
        splb_slv0_PLB_busLock: in     vl_logic;
        splb_slv0_PLB_RNW: in     vl_logic;
        splb_slv0_PLB_BE: in     vl_logic_vector;
        splb_slv0_PLB_MSize: in     vl_logic_vector(1 downto 0);
        splb_slv0_PLB_size: in     vl_logic_vector(3 downto 0);
        splb_slv0_PLB_type: in     vl_logic_vector(2 downto 0);
        splb_slv0_PLB_lockErr: in     vl_logic;
        splb_slv0_PLB_wrDBus: in     vl_logic_vector;
        splb_slv0_PLB_wrBurst: in     vl_logic;
        splb_slv0_PLB_rdBurst: in     vl_logic;
        splb_slv0_PLB_wrPendReq: in     vl_logic;
        splb_slv0_PLB_rdPendReq: in     vl_logic;
        splb_slv0_PLB_wrPendPri: in     vl_logic_vector(1 downto 0);
        splb_slv0_PLB_rdPendPri: in     vl_logic_vector(1 downto 0);
        splb_slv0_PLB_reqPri: in     vl_logic_vector(1 downto 0);
        splb_slv0_PLB_TAttribute: in     vl_logic_vector(15 downto 0);
        splb_slv0_Sl_addrAck: out    vl_logic;
        splb_slv0_Sl_SSize: out    vl_logic_vector(1 downto 0);
        splb_slv0_Sl_wait: out    vl_logic;
        splb_slv0_Sl_rearbitrate: out    vl_logic;
        splb_slv0_Sl_wrDAck: out    vl_logic;
        splb_slv0_Sl_wrComp: out    vl_logic;
        splb_slv0_Sl_wrBTerm: out    vl_logic;
        splb_slv0_Sl_rdDBus: out    vl_logic_vector;
        splb_slv0_Sl_rdWdAddr: out    vl_logic_vector(3 downto 0);
        splb_slv0_Sl_rdDAck: out    vl_logic;
        splb_slv0_Sl_rdComp: out    vl_logic;
        splb_slv0_Sl_rdBTerm: out    vl_logic;
        splb_slv0_Sl_MBusy: out    vl_logic_vector;
        splb_slv0_Sl_MWrErr: out    vl_logic_vector;
        splb_slv0_Sl_MRdErr: out    vl_logic_vector;
        splb_slv0_Sl_MIRQ: out    vl_logic_vector;
        aresetn         : in     vl_logic;
        aclk            : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of C_nfa_initials_buckets_REMOTE_DESTINATION_ADDRESS : constant is 1;
    attribute mti_svvh_generic_type of C_nfa_initials_buckets_AWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_nfa_initials_buckets_DWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_nfa_initials_buckets_NATIVE_DWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_nfa_finals_buckets_REMOTE_DESTINATION_ADDRESS : constant is 1;
    attribute mti_svvh_generic_type of C_nfa_finals_buckets_AWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_nfa_finals_buckets_DWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_nfa_finals_buckets_NATIVE_DWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_nfa_forward_buckets_REMOTE_DESTINATION_ADDRESS : constant is 1;
    attribute mti_svvh_generic_type of C_nfa_forward_buckets_AWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_nfa_forward_buckets_DWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_nfa_forward_buckets_NATIVE_DWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_sample_buffer_REMOTE_DESTINATION_ADDRESS : constant is 1;
    attribute mti_svvh_generic_type of C_sample_buffer_AWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_sample_buffer_DWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_sample_buffer_NATIVE_DWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_indices_REMOTE_DESTINATION_ADDRESS : constant is 1;
    attribute mti_svvh_generic_type of C_indices_AWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_indices_DWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_indices_NATIVE_DWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_SPLB_SLV0_BASEADDR : constant is 1;
    attribute mti_svvh_generic_type of C_SPLB_SLV0_HIGHADDR : constant is 1;
    attribute mti_svvh_generic_type of C_SPLB_SLV0_AWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_SPLB_SLV0_DWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_SPLB_SLV0_NUM_MASTERS : constant is 1;
    attribute mti_svvh_generic_type of C_SPLB_SLV0_MID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_SPLB_SLV0_NATIVE_DWIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_SPLB_SLV0_P2P : constant is 1;
    attribute mti_svvh_generic_type of C_SPLB_SLV0_SUPPORT_BURSTS : constant is 1;
    attribute mti_svvh_generic_type of C_SPLB_SLV0_SMALLEST_MASTER : constant is 1;
    attribute mti_svvh_generic_type of C_SPLB_SLV0_INCLUDE_DPHASE_TIMER : constant is 1;
    attribute mti_svvh_generic_type of RESET_ACTIVE_LOW : constant is 1;
end nfa_accept_samples_generic_hw_top;

library verilog;
use verilog.vl_types.all;
entity p_bsf32_hw is
    generic(
        ap_const_lv5_0  : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        ap_true         : vl_logic := Hi1;
        ap_const_lv1_0  : vl_logic := Hi0;
        ap_const_lv5_1  : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        ap_const_lv5_2  : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi0);
        ap_const_lv5_3  : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        ap_const_lv5_4  : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi0);
        ap_const_lv5_5  : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi1);
        ap_const_lv5_6  : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi0);
        ap_const_lv5_7  : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi1);
        ap_const_lv5_8  : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        ap_const_lv5_9  : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi1);
        ap_const_lv5_A  : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi0);
        ap_const_lv5_B  : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi1);
        ap_const_lv5_C  : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi0, Hi0);
        ap_const_lv5_D  : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi0, Hi1);
        ap_const_lv5_E  : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi0);
        ap_const_lv5_F  : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        ap_const_lv5_10 : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi0);
        ap_const_lv5_11 : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi1);
        ap_const_lv5_12 : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi1, Hi0);
        ap_const_lv5_13 : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi1, Hi1);
        ap_const_lv5_14 : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi0, Hi0);
        ap_const_lv5_15 : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi0, Hi1);
        ap_const_lv5_16 : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi1, Hi0);
        ap_const_lv5_17 : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi1, Hi1);
        ap_const_lv5_18 : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi0, Hi0, Hi0);
        ap_const_lv5_19 : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi0, Hi0, Hi1);
        ap_const_lv5_1A : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi0, Hi1, Hi0);
        ap_const_lv5_1B : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi0, Hi1, Hi1);
        ap_const_lv5_1C : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi0, Hi0);
        ap_const_lv5_1D : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi0, Hi1);
        ap_const_lv5_1E : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi1, Hi0);
        ap_const_lv5_1F : vl_logic_vector(0 to 4) := (Hi1, Hi1, Hi1, Hi1, Hi1);
        ap_const_lv32_1 : integer := 1;
        ap_const_lv32_2 : integer := 2;
        ap_const_lv32_3 : integer := 3;
        ap_const_lv32_4 : integer := 4;
        ap_const_lv32_5 : integer := 5;
        ap_const_lv32_6 : integer := 6;
        ap_const_lv32_7 : integer := 7;
        ap_const_lv32_8 : integer := 8;
        ap_const_lv32_9 : integer := 9;
        ap_const_lv32_A : integer := 10;
        ap_const_lv32_B : integer := 11;
        ap_const_lv32_C : integer := 12;
        ap_const_lv32_D : integer := 13;
        ap_const_lv32_E : integer := 14;
        ap_const_lv32_F : integer := 15;
        ap_const_lv32_10: integer := 16;
        ap_const_lv32_11: integer := 17;
        ap_const_lv32_12: integer := 18;
        ap_const_lv32_13: integer := 19;
        ap_const_lv32_14: integer := 20;
        ap_const_lv32_15: integer := 21;
        ap_const_lv32_16: integer := 22;
        ap_const_lv32_17: integer := 23;
        ap_const_lv32_18: integer := 24;
        ap_const_lv32_19: integer := 25;
        ap_const_lv32_1A: integer := 26;
        ap_const_lv32_1B: integer := 27;
        ap_const_lv32_1C: integer := 28;
        ap_const_lv32_1D: integer := 29;
        ap_const_lv32_1E: integer := 30;
        ap_const_logic_1: vl_logic := Hi1;
        ap_const_logic_0: vl_logic := Hi0
    );
    port(
        bus_r           : in     vl_logic_vector(31 downto 0);
        ap_return       : out    vl_logic_vector(4 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ap_const_lv5_0 : constant is 1;
    attribute mti_svvh_generic_type of ap_true : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv1_0 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_1 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_2 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_3 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_4 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_5 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_6 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_7 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_8 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_9 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_A : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_B : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_C : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_D : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_E : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_F : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_10 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_11 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_12 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_13 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_14 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_15 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_16 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_17 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_18 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_19 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_1A : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_1B : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_1C : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_1D : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_1E : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_1F : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_1 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_2 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_3 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_4 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_5 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_6 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_7 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_8 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_9 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_A : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_B : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_C : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_D : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_E : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_F : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_10 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_11 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_12 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_13 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_14 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_15 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_16 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_17 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_18 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_19 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_1A : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_1B : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_1C : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_1D : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_1E : constant is 1;
    attribute mti_svvh_generic_type of ap_const_logic_1 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_logic_0 : constant is 1;
end p_bsf32_hw;

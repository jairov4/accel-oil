library verilog;
use verilog.vl_types.all;
entity nfa_accept_samples_generic_hw is
    generic(
        ap_const_logic_1: vl_logic := Hi1;
        ap_const_logic_0: vl_logic := Hi0;
        ap_ST_st1_fsm_0 : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ap_ST_st2_fsm_1 : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        ap_ST_st3_fsm_2 : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        ap_ST_st4_fsm_3 : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        ap_ST_st5_fsm_4 : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        ap_ST_st6_fsm_5 : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        ap_ST_st7_fsm_6 : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        ap_ST_st8_fsm_7 : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        ap_ST_st9_fsm_8 : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        ap_ST_st10_fsm_9: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        ap_ST_st11_fsm_10: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        ap_ST_st12_fsm_11: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1);
        ap_ST_st13_fsm_12: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        ap_ST_st14_fsm_13: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1);
        ap_ST_st15_fsm_14: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0);
        ap_ST_st16_fsm_15: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1);
        ap_ST_st17_fsm_16: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        ap_ST_st18_fsm_17: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1);
        ap_ST_st19_fsm_18: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0);
        ap_ST_st20_fsm_19: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1);
        ap_ST_st21_fsm_20: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        ap_ST_st22_fsm_21: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        ap_ST_st23_fsm_22: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi0);
        ap_ST_st24_fsm_23: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        ap_ST_st25_fsm_24: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        ap_ST_st26_fsm_25: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi1);
        ap_ST_st27_fsm_26: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi0);
        ap_ST_st28_fsm_27: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi1);
        ap_ST_st29_fsm_28: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        ap_ST_st30_fsm_29: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi1);
        ap_ST_st31_fsm_30: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        ap_ST_st32_fsm_31: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi1);
        ap_ST_st33_fsm_32: vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        ap_ST_st34_fsm_33: vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        ap_ST_st35_fsm_34: vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi0);
        ap_ST_st36_fsm_35: vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        ap_ST_st37_fsm_36: vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        ap_const_lv1_0  : vl_logic := Hi0;
        ap_const_lv16_0 : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ap_const_lv64_0 : vl_logic_vector(0 to 63) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ap_const_lv1_1  : vl_logic := Hi1;
        ap_const_lv32_0 : integer := 0;
        ap_const_lv2_2  : vl_logic_vector(0 to 1) := (Hi1, Hi0);
        ap_const_lv32_1 : integer := 1;
        ap_const_lv64_1 : vl_logic_vector(0 to 63) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        ap_const_lv16_1 : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        ap_const_lv5_0  : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        ap_const_lv8_0  : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ap_true         : vl_logic := Hi1
    );
    port(
        ap_clk          : in     vl_logic;
        ap_rst          : in     vl_logic;
        ap_start        : in     vl_logic;
        ap_done         : out    vl_logic;
        ap_idle         : out    vl_logic;
        ap_ready        : out    vl_logic;
        nfa_initials_buckets_req_din: out    vl_logic;
        nfa_initials_buckets_req_full_n: in     vl_logic;
        nfa_initials_buckets_req_write: out    vl_logic;
        nfa_initials_buckets_rsp_empty_n: in     vl_logic;
        nfa_initials_buckets_rsp_read: out    vl_logic;
        nfa_initials_buckets_address: out    vl_logic_vector(31 downto 0);
        nfa_initials_buckets_datain: in     vl_logic_vector(31 downto 0);
        nfa_initials_buckets_dataout: out    vl_logic_vector(31 downto 0);
        nfa_initials_buckets_size: out    vl_logic_vector(31 downto 0);
        nfa_finals_buckets_req_din: out    vl_logic;
        nfa_finals_buckets_req_full_n: in     vl_logic;
        nfa_finals_buckets_req_write: out    vl_logic;
        nfa_finals_buckets_rsp_empty_n: in     vl_logic;
        nfa_finals_buckets_rsp_read: out    vl_logic;
        nfa_finals_buckets_address: out    vl_logic_vector(31 downto 0);
        nfa_finals_buckets_datain: in     vl_logic_vector(31 downto 0);
        nfa_finals_buckets_dataout: out    vl_logic_vector(31 downto 0);
        nfa_finals_buckets_size: out    vl_logic_vector(31 downto 0);
        nfa_forward_buckets_req_din: out    vl_logic;
        nfa_forward_buckets_req_full_n: in     vl_logic;
        nfa_forward_buckets_req_write: out    vl_logic;
        nfa_forward_buckets_rsp_empty_n: in     vl_logic;
        nfa_forward_buckets_rsp_read: out    vl_logic;
        nfa_forward_buckets_address: out    vl_logic_vector(31 downto 0);
        nfa_forward_buckets_datain: in     vl_logic_vector(31 downto 0);
        nfa_forward_buckets_dataout: out    vl_logic_vector(31 downto 0);
        nfa_forward_buckets_size: out    vl_logic_vector(31 downto 0);
        nfa_symbols     : in     vl_logic_vector(7 downto 0);
        sample_buffer_req_din: out    vl_logic;
        sample_buffer_req_full_n: in     vl_logic;
        sample_buffer_req_write: out    vl_logic;
        sample_buffer_rsp_empty_n: in     vl_logic;
        sample_buffer_rsp_read: out    vl_logic;
        sample_buffer_address: out    vl_logic_vector(31 downto 0);
        sample_buffer_datain: in     vl_logic_vector(7 downto 0);
        sample_buffer_dataout: out    vl_logic_vector(7 downto 0);
        sample_buffer_size: out    vl_logic_vector(31 downto 0);
        sample_buffer_length: in     vl_logic_vector(31 downto 0);
        sample_length   : in     vl_logic_vector(15 downto 0);
        indices_req_din : out    vl_logic;
        indices_req_full_n: in     vl_logic;
        indices_req_write: out    vl_logic;
        indices_rsp_empty_n: in     vl_logic;
        indices_rsp_read: out    vl_logic;
        indices_address : out    vl_logic_vector(31 downto 0);
        indices_datain  : in     vl_logic_vector(55 downto 0);
        indices_dataout : out    vl_logic_vector(55 downto 0);
        indices_size    : out    vl_logic_vector(31 downto 0);
        i_size          : in     vl_logic_vector(15 downto 0);
        begin_index     : in     vl_logic_vector(15 downto 0);
        begin_sample    : in     vl_logic_vector(15 downto 0);
        end_index       : in     vl_logic_vector(15 downto 0);
        end_sample      : in     vl_logic_vector(15 downto 0);
        stop_on_first   : in     vl_logic_vector(0 downto 0);
        accept          : in     vl_logic_vector(0 downto 0);
        ap_return       : out    vl_logic_vector(31 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ap_const_logic_1 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_logic_0 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st1_fsm_0 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st2_fsm_1 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st3_fsm_2 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st4_fsm_3 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st5_fsm_4 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st6_fsm_5 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st7_fsm_6 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st8_fsm_7 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st9_fsm_8 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st10_fsm_9 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st11_fsm_10 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st12_fsm_11 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st13_fsm_12 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st14_fsm_13 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st15_fsm_14 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st16_fsm_15 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st17_fsm_16 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st18_fsm_17 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st19_fsm_18 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st20_fsm_19 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st21_fsm_20 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st22_fsm_21 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st23_fsm_22 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st24_fsm_23 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st25_fsm_24 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st26_fsm_25 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st27_fsm_26 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st28_fsm_27 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st29_fsm_28 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st30_fsm_29 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st31_fsm_30 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st32_fsm_31 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st33_fsm_32 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st34_fsm_33 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st35_fsm_34 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st36_fsm_35 : constant is 1;
    attribute mti_svvh_generic_type of ap_ST_st37_fsm_36 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv1_0 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv16_0 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv64_0 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv1_1 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_0 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv2_2 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv32_1 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv64_1 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv16_1 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv5_0 : constant is 1;
    attribute mti_svvh_generic_type of ap_const_lv8_0 : constant is 1;
    attribute mti_svvh_generic_type of ap_true : constant is 1;
end nfa_accept_samples_generic_hw;

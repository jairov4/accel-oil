library verilog;
use verilog.vl_types.all;
entity system_nfa_accept_samples_generic_hw_top_0_wrapper is
    port(
        aclk            : in     vl_logic;
        aresetn         : in     vl_logic;
        indices_MPLB_Clk: in     vl_logic;
        indices_MPLB_Rst: in     vl_logic;
        indices_M_request: out    vl_logic;
        indices_M_priority: out    vl_logic_vector(0 to 1);
        indices_M_busLock: out    vl_logic;
        indices_M_RNW   : out    vl_logic;
        indices_M_BE    : out    vl_logic_vector(0 to 7);
        indices_M_MSize : out    vl_logic_vector(0 to 1);
        indices_M_size  : out    vl_logic_vector(0 to 3);
        indices_M_type  : out    vl_logic_vector(0 to 2);
        indices_M_TAttribute: out    vl_logic_vector(0 to 15);
        indices_M_lockErr: out    vl_logic;
        indices_M_abort : out    vl_logic;
        indices_M_UABus : out    vl_logic_vector(0 to 31);
        indices_M_ABus  : out    vl_logic_vector(0 to 31);
        indices_M_wrDBus: out    vl_logic_vector(0 to 63);
        indices_M_wrBurst: out    vl_logic;
        indices_M_rdBurst: out    vl_logic;
        indices_PLB_MAddrAck: in     vl_logic;
        indices_PLB_MSSize: in     vl_logic_vector(0 to 1);
        indices_PLB_MRearbitrate: in     vl_logic;
        indices_PLB_MTimeout: in     vl_logic;
        indices_PLB_MBusy: in     vl_logic;
        indices_PLB_MRdErr: in     vl_logic;
        indices_PLB_MWrErr: in     vl_logic;
        indices_PLB_MIRQ: in     vl_logic;
        indices_PLB_MRdDBus: in     vl_logic_vector(0 to 63);
        indices_PLB_MRdWdAddr: in     vl_logic_vector(0 to 3);
        indices_PLB_MRdDAck: in     vl_logic;
        indices_PLB_MRdBTerm: in     vl_logic;
        indices_PLB_MWrDAck: in     vl_logic;
        indices_PLB_MWrBTerm: in     vl_logic;
        nfa_finals_buckets_MPLB_Clk: in     vl_logic;
        nfa_finals_buckets_MPLB_Rst: in     vl_logic;
        nfa_finals_buckets_M_request: out    vl_logic;
        nfa_finals_buckets_M_priority: out    vl_logic_vector(0 to 1);
        nfa_finals_buckets_M_busLock: out    vl_logic;
        nfa_finals_buckets_M_RNW: out    vl_logic;
        nfa_finals_buckets_M_BE: out    vl_logic_vector(0 to 7);
        nfa_finals_buckets_M_MSize: out    vl_logic_vector(0 to 1);
        nfa_finals_buckets_M_size: out    vl_logic_vector(0 to 3);
        nfa_finals_buckets_M_type: out    vl_logic_vector(0 to 2);
        nfa_finals_buckets_M_TAttribute: out    vl_logic_vector(0 to 15);
        nfa_finals_buckets_M_lockErr: out    vl_logic;
        nfa_finals_buckets_M_abort: out    vl_logic;
        nfa_finals_buckets_M_UABus: out    vl_logic_vector(0 to 31);
        nfa_finals_buckets_M_ABus: out    vl_logic_vector(0 to 31);
        nfa_finals_buckets_M_wrDBus: out    vl_logic_vector(0 to 63);
        nfa_finals_buckets_M_wrBurst: out    vl_logic;
        nfa_finals_buckets_M_rdBurst: out    vl_logic;
        nfa_finals_buckets_PLB_MAddrAck: in     vl_logic;
        nfa_finals_buckets_PLB_MSSize: in     vl_logic_vector(0 to 1);
        nfa_finals_buckets_PLB_MRearbitrate: in     vl_logic;
        nfa_finals_buckets_PLB_MTimeout: in     vl_logic;
        nfa_finals_buckets_PLB_MBusy: in     vl_logic;
        nfa_finals_buckets_PLB_MRdErr: in     vl_logic;
        nfa_finals_buckets_PLB_MWrErr: in     vl_logic;
        nfa_finals_buckets_PLB_MIRQ: in     vl_logic;
        nfa_finals_buckets_PLB_MRdDBus: in     vl_logic_vector(0 to 63);
        nfa_finals_buckets_PLB_MRdWdAddr: in     vl_logic_vector(0 to 3);
        nfa_finals_buckets_PLB_MRdDAck: in     vl_logic;
        nfa_finals_buckets_PLB_MRdBTerm: in     vl_logic;
        nfa_finals_buckets_PLB_MWrDAck: in     vl_logic;
        nfa_finals_buckets_PLB_MWrBTerm: in     vl_logic;
        nfa_forward_buckets_MPLB_Clk: in     vl_logic;
        nfa_forward_buckets_MPLB_Rst: in     vl_logic;
        nfa_forward_buckets_M_request: out    vl_logic;
        nfa_forward_buckets_M_priority: out    vl_logic_vector(0 to 1);
        nfa_forward_buckets_M_busLock: out    vl_logic;
        nfa_forward_buckets_M_RNW: out    vl_logic;
        nfa_forward_buckets_M_BE: out    vl_logic_vector(0 to 7);
        nfa_forward_buckets_M_MSize: out    vl_logic_vector(0 to 1);
        nfa_forward_buckets_M_size: out    vl_logic_vector(0 to 3);
        nfa_forward_buckets_M_type: out    vl_logic_vector(0 to 2);
        nfa_forward_buckets_M_TAttribute: out    vl_logic_vector(0 to 15);
        nfa_forward_buckets_M_lockErr: out    vl_logic;
        nfa_forward_buckets_M_abort: out    vl_logic;
        nfa_forward_buckets_M_UABus: out    vl_logic_vector(0 to 31);
        nfa_forward_buckets_M_ABus: out    vl_logic_vector(0 to 31);
        nfa_forward_buckets_M_wrDBus: out    vl_logic_vector(0 to 63);
        nfa_forward_buckets_M_wrBurst: out    vl_logic;
        nfa_forward_buckets_M_rdBurst: out    vl_logic;
        nfa_forward_buckets_PLB_MAddrAck: in     vl_logic;
        nfa_forward_buckets_PLB_MSSize: in     vl_logic_vector(0 to 1);
        nfa_forward_buckets_PLB_MRearbitrate: in     vl_logic;
        nfa_forward_buckets_PLB_MTimeout: in     vl_logic;
        nfa_forward_buckets_PLB_MBusy: in     vl_logic;
        nfa_forward_buckets_PLB_MRdErr: in     vl_logic;
        nfa_forward_buckets_PLB_MWrErr: in     vl_logic;
        nfa_forward_buckets_PLB_MIRQ: in     vl_logic;
        nfa_forward_buckets_PLB_MRdDBus: in     vl_logic_vector(0 to 63);
        nfa_forward_buckets_PLB_MRdWdAddr: in     vl_logic_vector(0 to 3);
        nfa_forward_buckets_PLB_MRdDAck: in     vl_logic;
        nfa_forward_buckets_PLB_MRdBTerm: in     vl_logic;
        nfa_forward_buckets_PLB_MWrDAck: in     vl_logic;
        nfa_forward_buckets_PLB_MWrBTerm: in     vl_logic;
        nfa_initials_buckets_MPLB_Clk: in     vl_logic;
        nfa_initials_buckets_MPLB_Rst: in     vl_logic;
        nfa_initials_buckets_M_request: out    vl_logic;
        nfa_initials_buckets_M_priority: out    vl_logic_vector(0 to 1);
        nfa_initials_buckets_M_busLock: out    vl_logic;
        nfa_initials_buckets_M_RNW: out    vl_logic;
        nfa_initials_buckets_M_BE: out    vl_logic_vector(0 to 7);
        nfa_initials_buckets_M_MSize: out    vl_logic_vector(0 to 1);
        nfa_initials_buckets_M_size: out    vl_logic_vector(0 to 3);
        nfa_initials_buckets_M_type: out    vl_logic_vector(0 to 2);
        nfa_initials_buckets_M_TAttribute: out    vl_logic_vector(0 to 15);
        nfa_initials_buckets_M_lockErr: out    vl_logic;
        nfa_initials_buckets_M_abort: out    vl_logic;
        nfa_initials_buckets_M_UABus: out    vl_logic_vector(0 to 31);
        nfa_initials_buckets_M_ABus: out    vl_logic_vector(0 to 31);
        nfa_initials_buckets_M_wrDBus: out    vl_logic_vector(0 to 63);
        nfa_initials_buckets_M_wrBurst: out    vl_logic;
        nfa_initials_buckets_M_rdBurst: out    vl_logic;
        nfa_initials_buckets_PLB_MAddrAck: in     vl_logic;
        nfa_initials_buckets_PLB_MSSize: in     vl_logic_vector(0 to 1);
        nfa_initials_buckets_PLB_MRearbitrate: in     vl_logic;
        nfa_initials_buckets_PLB_MTimeout: in     vl_logic;
        nfa_initials_buckets_PLB_MBusy: in     vl_logic;
        nfa_initials_buckets_PLB_MRdErr: in     vl_logic;
        nfa_initials_buckets_PLB_MWrErr: in     vl_logic;
        nfa_initials_buckets_PLB_MIRQ: in     vl_logic;
        nfa_initials_buckets_PLB_MRdDBus: in     vl_logic_vector(0 to 63);
        nfa_initials_buckets_PLB_MRdWdAddr: in     vl_logic_vector(0 to 3);
        nfa_initials_buckets_PLB_MRdDAck: in     vl_logic;
        nfa_initials_buckets_PLB_MRdBTerm: in     vl_logic;
        nfa_initials_buckets_PLB_MWrDAck: in     vl_logic;
        nfa_initials_buckets_PLB_MWrBTerm: in     vl_logic;
        sample_buffer_MPLB_Clk: in     vl_logic;
        sample_buffer_MPLB_Rst: in     vl_logic;
        sample_buffer_M_request: out    vl_logic;
        sample_buffer_M_priority: out    vl_logic_vector(0 to 1);
        sample_buffer_M_busLock: out    vl_logic;
        sample_buffer_M_RNW: out    vl_logic;
        sample_buffer_M_BE: out    vl_logic_vector(0 to 7);
        sample_buffer_M_MSize: out    vl_logic_vector(0 to 1);
        sample_buffer_M_size: out    vl_logic_vector(0 to 3);
        sample_buffer_M_type: out    vl_logic_vector(0 to 2);
        sample_buffer_M_TAttribute: out    vl_logic_vector(0 to 15);
        sample_buffer_M_lockErr: out    vl_logic;
        sample_buffer_M_abort: out    vl_logic;
        sample_buffer_M_UABus: out    vl_logic_vector(0 to 31);
        sample_buffer_M_ABus: out    vl_logic_vector(0 to 31);
        sample_buffer_M_wrDBus: out    vl_logic_vector(0 to 63);
        sample_buffer_M_wrBurst: out    vl_logic;
        sample_buffer_M_rdBurst: out    vl_logic;
        sample_buffer_PLB_MAddrAck: in     vl_logic;
        sample_buffer_PLB_MSSize: in     vl_logic_vector(0 to 1);
        sample_buffer_PLB_MRearbitrate: in     vl_logic;
        sample_buffer_PLB_MTimeout: in     vl_logic;
        sample_buffer_PLB_MBusy: in     vl_logic;
        sample_buffer_PLB_MRdErr: in     vl_logic;
        sample_buffer_PLB_MWrErr: in     vl_logic;
        sample_buffer_PLB_MIRQ: in     vl_logic;
        sample_buffer_PLB_MRdDBus: in     vl_logic_vector(0 to 63);
        sample_buffer_PLB_MRdWdAddr: in     vl_logic_vector(0 to 3);
        sample_buffer_PLB_MRdDAck: in     vl_logic;
        sample_buffer_PLB_MRdBTerm: in     vl_logic;
        sample_buffer_PLB_MWrDAck: in     vl_logic;
        sample_buffer_PLB_MWrBTerm: in     vl_logic;
        splb_slv0_SPLB_Clk: in     vl_logic;
        splb_slv0_SPLB_Rst: in     vl_logic;
        splb_slv0_PLB_ABus: in     vl_logic_vector(0 to 31);
        splb_slv0_PLB_UABus: in     vl_logic_vector(0 to 31);
        splb_slv0_PLB_PAValid: in     vl_logic;
        splb_slv0_PLB_SAValid: in     vl_logic;
        splb_slv0_PLB_rdPrim: in     vl_logic;
        splb_slv0_PLB_wrPrim: in     vl_logic;
        splb_slv0_PLB_masterID: in     vl_logic_vector(0 to 2);
        splb_slv0_PLB_abort: in     vl_logic;
        splb_slv0_PLB_busLock: in     vl_logic;
        splb_slv0_PLB_RNW: in     vl_logic;
        splb_slv0_PLB_BE: in     vl_logic_vector(0 to 7);
        splb_slv0_PLB_MSize: in     vl_logic_vector(0 to 1);
        splb_slv0_PLB_size: in     vl_logic_vector(0 to 3);
        splb_slv0_PLB_type: in     vl_logic_vector(0 to 2);
        splb_slv0_PLB_lockErr: in     vl_logic;
        splb_slv0_PLB_wrDBus: in     vl_logic_vector(0 to 63);
        splb_slv0_PLB_wrBurst: in     vl_logic;
        splb_slv0_PLB_rdBurst: in     vl_logic;
        splb_slv0_PLB_wrPendReq: in     vl_logic;
        splb_slv0_PLB_rdPendReq: in     vl_logic;
        splb_slv0_PLB_wrPendPri: in     vl_logic_vector(0 to 1);
        splb_slv0_PLB_rdPendPri: in     vl_logic_vector(0 to 1);
        splb_slv0_PLB_reqPri: in     vl_logic_vector(0 to 1);
        splb_slv0_PLB_TAttribute: in     vl_logic_vector(0 to 15);
        splb_slv0_Sl_addrAck: out    vl_logic;
        splb_slv0_Sl_SSize: out    vl_logic_vector(0 to 1);
        splb_slv0_Sl_wait: out    vl_logic;
        splb_slv0_Sl_rearbitrate: out    vl_logic;
        splb_slv0_Sl_wrDAck: out    vl_logic;
        splb_slv0_Sl_wrComp: out    vl_logic;
        splb_slv0_Sl_wrBTerm: out    vl_logic;
        splb_slv0_Sl_rdDBus: out    vl_logic_vector(0 to 63);
        splb_slv0_Sl_rdWdAddr: out    vl_logic_vector(0 to 3);
        splb_slv0_Sl_rdDAck: out    vl_logic;
        splb_slv0_Sl_rdComp: out    vl_logic;
        splb_slv0_Sl_rdBTerm: out    vl_logic;
        splb_slv0_Sl_MBusy: out    vl_logic_vector(0 to 6);
        splb_slv0_Sl_MWrErr: out    vl_logic_vector(0 to 6);
        splb_slv0_Sl_MRdErr: out    vl_logic_vector(0 to 6);
        splb_slv0_Sl_MIRQ: out    vl_logic_vector(0 to 6)
    );
end system_nfa_accept_samples_generic_hw_top_0_wrapper;
